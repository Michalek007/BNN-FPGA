-------------------------------------------------------------------------------
--
-- Title       : layer_hidden
-- Design      : uart
-- Author      : Michal
-- Company     : AGH
--
-------------------------------------------------------------------------------
--
-- File        : C:\Users\Public\Projects\MyDesigns\uart\src\layer_hidden.vhd
-- Generated   : Tue Feb 13 20:33:23 2024
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {layer_hidden} architecture {layer_hidden}}

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.numeric_std.all;
use work.layer_constants.all;

entity layer_hidden is
	 generic (
		 N_INPUTS : integer := LAYER_HIDDEN_N_INPUTS;
		 N_OUTPUTS : integer := LAYER_HIDDEN_N_OUTPUTS;
		 POP_CNT_MAX : integer := LAYER_HIDDEN_POP_CNT_MAX
		);
	 port(
		 INPUT : in STD_LOGIC_VECTOR(0 to N_INPUTS);
		 OUTPUT : out STD_LOGIC_VECTOR(0 to N_OUTPUTS)
	     );
end layer_hidden;

--}} End of automatically maintained section

architecture layer_hidden of layer_hidden is

component pop_cnt
	generic (
		N_INPUTS : integer := N_INPUTS;
		N_OUTPUTS : integer := POP_CNT_MAX
	); 
	port(
		INPUT: in STD_LOGIC_VECTOR(0 to N_INPUTS);
		OUTPUT: out STD_LOGIC_VECTOR(0 to N_OUTPUTS)
	);
end component;


type WEIGHTS_ARRAY is array (0 to N_OUTPUTS) of STD_LOGIC_VECTOR(0 to N_INPUTS);
type POP_CNT_ARRAY is array (0 to N_OUTPUTS) of STD_LOGIC_VECTOR(0 to POP_CNT_MAX);
type NORMALIZATION_ARRAY is array (0 to N_OUTPUTS) of INTEGER;

signal W: WEIGHTS_ARRAY;
signal W_XOR_INPUT : WEIGHTS_ARRAY := (others => (others => '0')); 
signal POP_COUNTER : POP_CNT_ARRAY := (others => (others => '0'));

signal GAMMA : NORMALIZATION_ARRAY := (25, 287, 8, 260, 923, 291, -20, 286, 609, 1340, 250, 955, 8, 0, 1169, 910, 28, 1289, -4, -11, 36, 25, 18, 182, 366, 141, -18, 570, 864, -20, 10, 5, 206, 1028, 1060, 11, 343, 286, 2, 23, 9, 116, 9, 1095, 117, 792, -7, 0, 9, 155);
signal BETA : NORMALIZATION_ARRAY := (-5, -5, 2, 4, 111, 4, -3, -3, 79, -144, -1, -54, 9, 0, 64, -119, 3, 92, -1, 0, 5, 0, 6, -3, -102, -7, -5, -16, -40, -6, 0, 0, 4, -91, 52, 0, -6, -1, -9, 9, 0, -14, 0, -65, -7, 4, 0, 0, 3, 29);
signal MEAN : NORMALIZATION_ARRAY := (0, 0, 0, 0, 12, 0, 0, 0, 7, 7, 0, 7, 0, 12, 8, 11, 0, 9, 0, 0, 0, 0, 0, 0, 13, 0, 0, 14, 10, 0, 0, 0, 0, 7, 12, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 9, 0, 13, 0, 0);
signal STD_DEV : NORMALIZATION_ARRAY := (1, 1, 1, 1, 54, 1, 1, 1, 48, 69, 1, 56, 1, 59, 49, 66, 1, 66, 1, 1, 1, 1, 1, 1, 41, 1, 1, 52, 66, 1, 1, 1, 1, 44, 64, 1, 1, 1, 1, 1, 1, 1, 1, 57, 1, 54, 1, 53, 1, 1);

signal NORMALIZED_BATCH: NORMALIZATION_ARRAY := (others => 0);

begin
	
--	--	simulation
--	W(0) <= "00000000";
--	W(1) <= "00000000";
--	W(2) <= "00000000";
--	W(3) <= "00000000";
--	W(4) <= "00000000";
--	W(5) <= "00000000";
--	W(6) <= "00000000"; 
--	W(7) <= "00000000";

	
W(0)<="11011101101001101011111111101111110011010011111110";
W(1)<="11111010001011101011110111111110100011110011111110";
W(2)<="01011101101111111011011001111111110111010111101110";
W(3)<="00101011101111111111111111111010110110010101111011";
W(4)<="00001001110100011110101000001010001100111001100001";
W(5)<="00111000000000101111011101111111110111010001111110";
W(6)<="11101110101010111011110111110110111011110111111110";
W(7)<="11101000101101111111011100111101010011010111111110";
W(8)<="01011100111001010010101001000110000100111010110011";
W(9)<="10001110011000111010011011010010100000101011010000";
W(10)<="11111011101100110011010101010111110011110011011110";
W(11)<="11101010111010100110100111100001000001001110000110";
W(12)<="01100110101111110011111000111100110011110110101111";
W(13)<="00110010011000010000100111000100100000101010010010";
W(14)<="10110100010100010100011110001011101100101100011001";
W(15)<="11000011010100111000101101100001101000001001110000";
W(16)<="01111001101111110011011100111111110111010001011110";
W(17)<="00001111010011111100001111110010100000111110010100";
W(18)<="11100111101111011011011101110011111111010010011110";
W(19)<="11011011001010111011110110111111110111110100111101";
W(20)<="11011111101011101001011011110011110111010101111111";
W(21)<="11111001001010111011011111111111111111010100011110";
W(22)<="11101100001001111011010110011111011111110111111111";
W(23)<="11111111001110101001110111111111011011111111111110";
W(24)<="10101000110110110100011111001000000000001000011001";
W(25)<="01111110101110111011111001111111010011110111111111";
W(26)<="10011100101101111011011111111111111110010111101101";
W(27)<="11101011010011010110100101000010100100101000000001";
W(28)<="01110000111000000000100111100001100000101100010010";
W(29)<="11111110001011111111011011111110111111100010101110";
W(30)<="11111111001110111011010001010111111111110111111111";
W(31)<="11011101001111101111111001110110010011010111111111";
W(32)<="11011000100111111011011011111110110111110111111101";
W(33)<="00011100111010010010000010011101000000111011110011";
W(34)<="10011011011110000110000010001001000001011010100001";
W(35)<="01011011001101101011111101111101110111010011011111";
W(36)<="11111100001100101001111110111101110111110011111010";
W(37)<="11101111001111111011110101111110110011110011111110";
W(38)<="11011000001100001011110111110101010111110011111010";
W(39)<="01111101101010111111111111111101011111110101011110";
W(40)<="11110101101000101111111111011111110011010110111111";
W(41)<="01011111101100111011111100111101010111010111111110";
W(42)<="01101110000111111111111111011111111111110111111110";
W(43)<="10101010011100110111100111001001000000000000100000";
W(44)<="01111110101101101111011110011111011111000111111101";
W(45)<="10011100110010010100001110011100000001011110010000";
W(46)<="01111110101110101011111110111111110110110110011010";
W(47)<="10111000110111010100001110001001001001001100010001";
W(48)<="01110011101110111111111110111111111011110010111100";
W(49)<="01100000101111101011110000110111010111110001101110";

	W_XOR_INPUT_i:
	for i in 0 to N_OUTPUTS generate  
	begin
		W_XOR_INPUT(i) <= not (W(i) xor INPUT);
	end generate;

	POP_CNT_i:
	for i in 0 to N_OUTPUTS generate
	begin
		pc: pop_cnt port map (INPUT=>W_XOR_INPUT(i), OUTPUT=>POP_COUNTER(i));
	end generate;

	NORMALIZED_BATCH_i:
	for i in 0 to N_OUTPUTS generate
	begin
		NORMALIZED_BATCH(i) <= GAMMA(i) * (to_integer(unsigned(POP_COUNTER(i))) - MEAN(i)) / STD_DEV(i) + BETA(i);
	end generate;
	
	OUTPUT_i:
	for i in 0 to N_OUTPUTS generate  
	begin
		OUTPUT(i) <= '1' when (NORMALIZED_BATCH(i) > 0) else '0';
	end generate;

end layer_hidden;
