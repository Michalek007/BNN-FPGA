-------------------------------------------------------------------------------
--
-- Title       : layer
-- Design      : uart
-- Author      : Michal
-- Company     : AGH
--
-------------------------------------------------------------------------------
--
-- File        : C:\Users\Public\Projects\MyDesigns\uart\src\layer.vhd
-- Generated   : Wed Feb  7 03:50:28 2024
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {layer_input} architecture {layer_input}}
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use IEEE.numeric_std.all;
use work.layer_constants.all;


entity layer is
	generic (
		 N_INPUTS : integer := LAYER_INPUT_N_INPUTS;
		 N_OUTPUTS : integer := LAYER_HIDDEN_N_INPUTS
		);
	port(
		INPUT: in INPUT_ARRAY;
		OUTPUT: out STD_LOGIC_VECTOR(0 to N_OUTPUTS)		
	);
end layer;

--}} End of automatically maintained section

architecture layer of layer is

type INTEGER_INPUT_ARRAY is array (0 to N_INPUTS) of INTEGER;
type INTEGER_W_DOT_INPUT_ARRAY is array (0 to N_OUTPUTS) of INTEGER_INPUT_ARRAY;

function f_sum (x : INTEGER_INPUT_ARRAY) return integer is
   variable n : integer;
   variable sum : integer;
   begin
      n := 0;
	  sum := 0;
      while (n < N_INPUTS+1) loop
		 sum := sum + x(n);
         n := n + 1;
      end loop;
      return sum;
end function;

type WEIGHTS_ARRAY is array (0 to N_OUTPUTS) of STD_LOGIC_VECTOR(0 to N_INPUTS);
type W_DOT_INPUT_ARRAY is array (0 to N_OUTPUTS) of INTEGER;
type NORMALIZATION_ARRAY is array (0 to N_OUTPUTS) of INTEGER;

signal INTEGER_INPUT : INTEGER_INPUT_ARRAY;
signal INTEGER_W_DOT_INPUT : INTEGER_W_DOT_INPUT_ARRAY;  

-- weitghs
signal W: WEIGHTS_ARRAY;

-- dot product of weights and input
signal W_DOT_INPUT : W_DOT_INPUT_ARRAY := (others => 0);

-- dot product after reLU activation function
signal RELU : W_DOT_INPUT_ARRAY := (others => 0);


-- normalization params
signal GAMMA : NORMALIZATION_ARRAY := (389, 1683, 973, 966, 1194, 724, 1227, 958, 1030, 1089, 787, 772, 1431, 1011, 490, 1266, 984, 1233, 389, 1128, 867, 1321, 1350, 932, 792, 458, 935, 1132, 1035, 854, 1207, 1287, 835, 1486, 1200, 1427, 1144, 1540, 1704, 1342, 796, 1096, 988, 953, 956, 1462, 1303, 1254, 1075, 785);
signal BETA : NORMALIZATION_ARRAY := (212, 78, -567, -1034, -434, -443, -446, -513, -398, 1035, -600, -17, -533, -1063, -472, 82, -1002, -201, -319, -585, -657, -501, -456, -618, -265, 66, -333, -113, -1000, -458, -1008, -569, 415, -737, 271, -543, -178, -195, 217, -381, 1158, 78, -16, -146, -386, -289, 67, -247, -715, -10);
signal MEAN : NORMALIZATION_ARRAY := (851, 1630, 1420, 0, 1051, 2029, 1201, 603, 1008, 0, 1448, 2299, 641, 0, 4351, 4918, 0, 1914, 3221, 359, 1152, 1107, 594, 1654, 1963, 185, 2233, 1851, 0, 3457, 0, 726, 9348, 417, 4110, 917, 1966, 1804, 2722, 812, 0, 2510, 2691, 2494, 1995, 1701, 2192, 1848, 191, 3735);
signal STD_DEV : NORMALIZATION_ARRAY := (2860884, 7092279, 4950837, 1, 4161015, 5325279, 4045026, 1699480, 4581017, 1, 5379040, 8057932, 2881993, 1, 9718124, 17176330, 1, 5906370, 9058869, 972429, 3469561, 4369966, 1610694, 4992200, 5516197, 791325, 7131961, 5685812, 1, 8836900, 1, 3309160, 14098976, 1183727, 11977026, 3394908, 7312852, 7162826, 10895340, 2952647, 1, 10902672, 8625509, 5510024, 6202531, 6572673, 8599154, 7533063, 465358, 13204256);

-- normalized relu
signal NORMALIZED_BATCH: NORMALIZATION_ARRAY := (others => 0);

begin

--	--	simulation
--	W(0) <= "110";
--	W(1) <= "110";
--	W(2) <= "110";
--	W(3) <= "110";
--	W(4) <= "110";
--	W(5) <= "110";
--	W(6) <= "110"; 
--	W(7) <= "110";

W(0)<="0011010001101101001110010011111111111111111001111111010001111111111111110101111000110101111110110010101111111010011110000010001010111111110110110000000011111111111011000010000001100000000110011110000000101010000000111111101101000001001100000111001110111110010000000000111100011110111000000010001111110001111111110000000100111100001111111000000000111011100000010110111000000111100000001000001011110011111111100001000110001111111111111100011000110000100111111110110000010010000110000111110111000000010010010000001110011100010000001000110000111001100000000001101111000011000111000000000110101110011101100011111111111001110000101001111111111111111000000001100111111111111110100010001101111111111111110110100111111111111110001111100100111000110111000100111000000111111101110100101110111101";
W(1)<="0000100101111111111111010110101001001011111111111111001010000100111111111111111111100111111100111010001111111010111111001110000111111111110101111111111111111111111100000101111111111111111111111001001111111011111100111111100001011110011011000000011110100111101010100000000000111011101110001100000000000001111100011111100000000000001010010100001100000000000011111001010000011000000000111011110010000000010000000010100111101110000001000000011100001111111000000100000001000000111111110000001100001000010011111111100101111111100000011111111111111111111111100111111111111110011101011111111111111111111111101001011111111101111111111101011111011111011111110000111111111111111110000000000010011111111111101011110000000000000011110100101111010010011110010101001010101001001110100100001110110010";
W(2)<="1001111111110111111111110011110111111110011110111111010100001111100000000011111111001111000000000100001000100111110000000000000000000000111001100000000111011100000010101100000011111111010000000001100000000111111111000000001010010010011101111101010011011011011001111111110110100110101010100010011011001000001000000100010001010110000011100011111111011100000001001011111111111111110000010000110111111011101101100111111111111011101001111111111111111110000111101001111111111111111001001000000011110001111111110000000000001110000001110111100000000000000000000011111100000000000000000000001111100000000000001100101000110101100000000011100101110101011100001111111111100111111111111011111111111111011101101000001111101011111111111111110111101100111111111011111110011010100001010111000011101010";
W(3)<="0010000011110110001011010011100001000111011011011100011010100100011100100100000111010010111111110100000011100110101111100011000111111010011101011111000000000010101101010111111101000000110011011110111101100000001000000100001100110100101100100000000000110100010000110000000100000100111101000110100010000110100110100111101000001000010001111100011100000000010000011001110011001000010000000011110010000100110010000000001111001010100111110001100000111101010100001011101100100111000011011110011000100000000001010111010111001000000000100001110001000010101000000010101111100000011110010000101111111010000100011011100011111111000001100000010110111111101111000110010000000110110000011110001101101000000110011111011001111001011001100111000101100111101000001110100010101011111001001111101101101101";
W(4)<="1000111111101111000000000110111111111111111111111111101010011111111101111011111110111000000000000000000111111110000110000000000000000011000000111000000000000000000000110011000000000000000000000011010100000000001000000000010011000000000000010000000001011000000100100101100000000111100000011001111010110011010100000111011100000100110111010000011111111000010101001011001011011001100001100111011000000010111110000000101111100000011111111000001011111110100001111111111011111100110010000111111111111100011111101000000110101111111101111010000000010111111110111100001010010000111111111101100111101100001001111111011111001101010000000000000000000000000001111000000000000000000010000010000000000000000000111001100000000000000000000011001010000000000000000000000100001100000101011110110000111110";
W(5)<="1100000110111110111110001011001000000001000101000000000001100000000111000000000001000111011111111111100000000101111111111101111110010000000100111111110001111111111110110111110110101001111111001011111110011000110111111100001001111010011011111111110000110111110111000111111110000000111110000111011111100000000111100000000011110100000000011110000001000111100000000000110000000010011000000000010011100000000000100000000001111111000010100100000000010111111100001000001111111111000111111011101111111111111000010111110011110011101110100011111111111000001111100010011111111110100000111001011000111001111010000011000110100010111000100010101110101100011110000000000001111110000001001100100000000000011110000100100000000000000000010001001100000000000110000000000001011010111001111100011010111010";
W(6)<="0100000100001000000101100011100100000000000000000000011111100000000000000000000001101111111100100101000000000000011101111001000100000100001001110111111000000011111110100111101011000001111011111011111110011101010010000111101011111000000011100011111100111111010100100111000011111010111110010000111101111111111111111111000011111111111110011111000000011111101111111100011001000100111100100000000101110001001001000000000001110110000001011100000000000111100000001111100000000000100010000000010110000000000001111000010001011100000000100110100000011110111101100000001100000001110111110000000000110000011101011111100010000011100000100111011111101010011010000000001101111111111001100100000000000011111110101000001100000001101100110101110010100000001111000000111111110100101111010001111001001110";
W(7)<="1110111111111111111110110101010000001110100000010010011100100000000110000100001110101110000000110111111011100001001000010100101001101100000101100000000010100111000000000000000000101000111100000110010000000000010001000000011000000000000000100000110001111110000001110110000010010101011111001111111000001011010000000111111111000001110100010011111111111000000011111101001111111101100001111011011001111100001100000110011101110001111001110000100111011110100011101111000110100111111000000111011100010110101111100000010111110001100101111110000011000010000111111111111000001010010000011111111111100000111110000001111111111111100011110110000011111111110011111111001001100010111110000111110000000001110011100010110001110010000100000011101001100000000000000000001111000001101100100000001001001100";
W(8)<="0000111110100000000111110101010111111111111111111110010100100011111111010001111110011100000010101101011101111010100000001111111111110001001111000000010111110010011000000100000001011111110001100001000000000000111111010110001110000000101000011101000001000000111010110000011100000100011111000010000001110010000110001110101000000011100000010011111100100000001010100001011111010000000001110010010100011100000000001111011101111001111111100001111111111110000111111100011111111111110100000011111111111111111111101000001000111111010111111110000001000010000000001111111000000011100000000000011111100000001001000100000000101110100000100101111101010000111000101001101010110111111110111011110111111111111111111101010111111111111111111110101010001111111111111111110000111111111101101110111101000101";
W(9)<="1011001010100000001101010010000111011010100100111111011100101100110010110101100010010110101010011111001001011000011000010111000111111110100111111101000010110010101000111100000111001010110001010111101001010011000010001011111010100000001101001101100000100010100000000010000001000000111100001100011000010101100000010100100100001100010111011100101110110100011011101011100000001000100010110110111110101100011001010001010111101001000010000101001001000110111011100100001010110110000001010000111100000010000010101001100000011001111101001100001011010000010000110001110100010010011001111000100010010000100000100101000101000000001110010000000001001001001100010011010000011000010111010100111001110000101011111100111100111111011100010000111011101001001010010011010011111001001001010001010011100100";
W(10)<="1100100100000000110110100100010100000000000000000000011010100000000000000000000001011010000000000000000000000001011000000000000000000000011011100000000010000110100111001111111110011000010100011110111111111101111011011111111001111111111111001011101100110111111011111111110110110000111111110111111110111111010011111100111111111110101110001111100010101111111111111001111110001000111111001000000011110001100011100000000001101000001110010000000000000110000000010000000000000000000000000001000100001000000000010000000100011000010000000010000000000011111001100100011111000000001110000010111001101110011000111000010000101101010000111011100011010100111000000010110010011111110001111011111000010010011000001010001111000101011100011101110000111111100111010000111010101100011000000011000111110111";
W(11)<="1111000011101111000001110110000111111111111111110011101010011111111111111111111111110111111110001010111011111101011111011100101000001111111010010000111010000101111111001010100010111000001001111110111110011101010000111101100011101011111111000001101110001110011111111100000000011110111111101111110000000001111111111110111100010000000111111111001100111100000000011010011000001111011000110001101011100000011111101110000110000110000111111111000000011100100000011111110000000000110010000001111111000000011110000000000101111100000111111010000000001111111001001111101010000000101011110001011110100000000001001110111111111000000000000000001111011111110010000000111101111111101111111010000001111111100000111100101000000101100000000001010111001000010001000000001111000010001111100000011011101110";
W(12)<="1101110000111000111111110101001000000000010001000000010001000010000000000000010011011000000000000000000000010010010000000000000000000100101111000000000000000000000010101110000001111111100000000001110011110000111111100000000101111111111111011111100000101011111111110111111110000100101111111111001011100110010011111111111011001100010001111011010101101110110100100010111111110101111111101100010111111010011101111000000001011001101000110000000100010001000110101000010000000011010100010111110001001011000100010001001100000100000000000100001000000000001001000000010111100000000000010100000101111111000000000000001100000000011000000001000000110011000100000001110010001100100111001011111111111110111101011011101111111101111111111000100111101101101110011001111110101101111100000000100111000100";
W(13)<="1110111110100000000011010001011010101111001000100100010000000011011000010000111110110111110010101101010011000110000010001100101110111010010010100010100000011100011110100100100100000000000000000101100000100010010011000100101001010000000010100100001011011111011000000000110100001110110110110111100110011000100000011111110000000001001011110001101100000000101001001100010011000010000000000000110111110010000001000000000001000101110000011110010100001100110111000000001101000010011101000000001100101101000110010111101110000000001010111100111110100101000000010110010001101011001111000011111000011110100010001110011111000000110101100011110101111011100000111010110000000111001011011101110110000010011100110101010110110110010100000101110100111100000101000110100101010010111010000101100010011011";
W(14)<="1110000000101110110110001011000000000010000000000000100101100101100000000111110001011111111000011111101111011110011111111111001000100111110001110111111010000110110111000111111011111010010011011110111011111111100000111111111001111110011110000111001110000111111111111010000001111110111111111110011100000011111011111111111111111010000111101111000010011111100000011100011000000101111110100000001010000000111111110000000010101010000111101111000000000011101000011110111100000011001100000111111111000000011010000100111111110100001010010001111001111100001111100001101111100000110110010000001110111110000101011011110000011010111000011011001100011111110010000000010111111111111110111100111111111111101101111111000110011111110100000000011101001000111111000000001010010111101100100100100000011010";
W(15)<="1000100010011100100000110001101010000111001000000000111111100000110111111100000000110111010011111111001100001100011111111111111110100111110011111111111111100110111111100001111111111111011111011111000111111111001111111110110001011111011110111111111111000100110000010111010111111110100000000010001110000011111001000000000011111010000111101000000010001111100000001111110000000111111100000000000111100001010111100000000010011111100000001110000000110001111111001100110000000011000011111100001100000000111100010111111110110000001110010001111111110101010111001111100011111011010111100101101010001111001111011101111111101000111101111111111110111100100010010000010111111111100001001000011111111111000000110110010000000111110110000000001000001000001111110001011001001111001000011111110101111101";
W(16)<="1010000010100111010001111100000101100101111000101001010000011011111100111010110001111010110101111000010101100011011101010010000101100110111101000110001100110000000010110111100011000011000011101000100001100110101110010111111011000010000000000010011110000101000011110000001000011011011000100100110110110110101001001000000001000110001001111110011001111100100001110011011101100000000001000111110010001010101101100000001111101001000110000011100100010110001101001000101000101111101101100001000100001110010001100111001000010001000110000001000110110010000000011111010111000110000010100001000010010100110100101000001100010010000010000101000110101011010110101110011000010100000101000001000000100101001001100011001000000100110000101110111011011110000111110000100010000010000100011000101001000000";
W(17)<="1101111111111011001100011011100101111111111111111110000010000010100100111111111110010110000000000000011111111110010000000000110111111010010111100000000011100111101000001110000000000111010000110101010000000001010000100000111100000000011111100000100111101100000001111110000010011111110000001110011000001110111110000001111101010000101110111000000011101111100010000011011000000000011000000111011000000000000001100000001111101100000001111110000010111111111110101111111000000011111011111111111111100000001111110111111111111111000101111110110111111111111010011000001001111111111110010110100111111001001110000011101000011101100100010000000001000001011101111111100111001000001111000101111111100001000000111100011111111101100000111101001101010111110011011110101001111101011011000110110101101100";
W(18)<="1001100111100010010001110101111100011000000110000000000011100000111110001000000001011111000011111111000000000001101011100011111110100000000101001110000111111011110001010111111100000010101111100111001111111010111111111011000001111111111011111111001000011111110111101011100001100000111110000100000110000110000111000000000000100011000000001101100000000010011100000001110000000000001111000000010111100000110000011111001001111111101111000011111111101110111100101000001111111110000011111111111000111111111111010111111001110011111111100001111111111111001110111000010110111110111000111011100000001011110011000011110110000000011001111111011110111000000110110000010010001000000001101000000000000000001000001000000000000000000000001100100111010000001110000010010110001001111110101000001000000100";
W(19)<="1000000000010100000010001001101111111110000000000000010011110111110000110111111100100110000110110110111111111101100100101111000110101011100010000001011110000111110111000000000001100000110000011110100000110101010000000101110010100011111100000000001111101000111100110000000100101101000111001000000000001001011000011111010000000000000111110011111100000110101000010101101100100000011100100001101001100000000011110111000010100010000000011111100000001001010000000011111100000000111101000000111111100000001011010000000001111110000000111000100000001111110001001111100010000000000000010111101110100000000011010011010101111110000000001101101011111111101111000000111111111111111111101100000000111111110111111100101011111001111100000000000111000011100111110011000111100010101001111100100001001010";
W(20)<="1101100111111111110011111101001100001111110111111111001001100000000111111111111111001111001000001110011111110101011001111100000110001111001011101001110011111111101101101111110011110010101001111101111110000010001110101111111001110010000001111111011110110111000001010011111110110000111100100111111101111111000111111000001001110110000000011111010001000011110000000000111100000000000000000000010011110000000100000000000001111010000001100000000000000110000000101010000000000011011110000011011000001111111100101000010001011111111111111010000001110010111111111111111000000111101111111111111001101000000000011101110111100010010001010110011111111101011010000011100010111111100001001110011001000011111100101011010110010110000110110001011000100011111111100000010010001000101111011111001110000010";
W(21)<="0100111100011011111101110001011010000000000000000000111011100000000000000000000000100110000000000011011000000011111000000010011111000000001001100010010000001110111101100111011101001000011111010110111111111000100001111010001111111010000011001111110100111111100110000000111110110001111101110001100011111010010111111010100010011111111000011111100010000001111110110010111111000100011110001110001111111111000100000000000001111111111111000000000000000010100111111100001000000000000100001111111000111001000000010000110111100110111000001000000011101111110101000000110011001110111101000100000101001000001011111111000000001000110000010111111100000000101000000000001111111000110011011110000000111111111110001010100110000001001110011100110110111000001110001011110010111001010110010000001000011110";
W(22)<="0100100110011111010100000111111000000001110111111000001111100000001111011111001110111111000000000100010011110011001000000000010000001111000010110111000011000100011101010011100110111111111101111101101100111010011111100001010010111111000000111111000101001111000000000111101100000011011100000001001101111000001000000000001111101010000000100100001001010100000000000001011000101101000000000000011001100000001000000000000001101000000000010000000000011100000000000001100000001110010110000011111111000011010001101000001001111100111111101110100000011011110001011011111110000111101101001111110011001000010000011110011111100011100001110100110000111110000011001011101111100111100000101011110010111100011110000100011111111111111111001100001011101011111111000001000000010110000111100000010110001100";
W(23)<="1010111111111111111111100010000111111111111111111111010111110111111111111111111110000100000011101110111111101001000000011111111101000011000000000111111011111001100100110000111111111110010111110011100111011111010000000000010010011110010011000000000101011001101100101100000000001010000010100111110000000000100000000110110011000000000010001000001101110110011000001101000000010110010001100111010111000000010001001110011111111100000000000001111111111110111000000000011111001111110011100000000001111110100111101111000000000111100000001110011111011100111111111001110011111111100001111100110111001111110001001110001001110100111111110000110111110110000100101110110111111000010000001001111111111110000000110111101111111111111110000000101011011101111111111111111001001100000000001100101101001100";
W(24)<="1011000000000000000000000001100000010000011001111101001100011101011111001111000000110000111111001001111110000101100011111111000101010000010010001101011100100100000100011001101110011000000000000001000111101111100000000010010110010000100111000000011100011000000110111100001000100001000000001101110010111000000000001101111110011001100000000000111011111000100101011110000001111111100010011111101100000111111110011101111100000000000011111011111111110000010000000001000111111111000001000000000000011110100000000010000000000001100000000001011100000101001110110000000101111111111111101100000001100111111110100101101000000111011111110110000111100010001011111111111100011100111100000110111111100000000011100000101011111111011010110111100110000111000000000011100101001100011101111110001100100110";
W(25)<="0000111111111111110001111110010011111111111111111111101011111111110011001111111110111100101000001000011100111000100110000000100001000000011010010000000000010111111001010100000000000001010000110001100001000000000101100010001100000000000000000010101001110000001100000000001111110101100011100000000000011111010100001101000000000001111001010001101000000000000111100010101110100000000000011110010010001100000000000011111111110001111100100000000101111100000111111110000001011100110000001111111111100010010111001000110111111110000111111110100011010111111101111111101000000111111111011100111111100000011011110010110001011100010000111011111111001001111101100010100011111101000110110000000000111100000000000000110001000000000000000110001001000111111110111000011011101011011100011011011001100011";
W(26)<="0110111111100100110000111100100111111111111111111111101110011111111111111111101011011000111111111111111100000010000111011000000000000000000011011000000111110000000000001100000101111111010000000010100000111100111101000000100110000000101101011101000011110000010111010001111110000101000001001100000111111100010000001101000010011000010000100001101100000001110011000010000111110100100011111110000000011111010110001101111100000001111101110001011011110000000111111100001011111110001101000000000001100101110000111000000000001111111111000010000000000001111111010100001100000000001111111110100000100000000001111110101000000101000000111100000000010000010111001111111111000101010010000111111111111111111111111001011111111111111111111110110101001111111111111111110111001011101100101011001000000110";
W(27)<="1000111111101100000000000100110111111111111111111110100010011111111111111111111100111000111111111110011110000000100111100011111000011000000110011000000001010001000000001001000100000000000000000000011100001000000001000000010111000000101001100110000001000000000001101110111000000111000000000100000111000000000100000000001100110000001111010000000000010110000000011010000000000001111000010101000000000111111111000011111111010000111111101100011111111011100111111110111001111111001010000110100111111001111001011000000001111111011111001111100000000111111101000011101010000011011111111100000111011000000011111111100000000001010101100000101000000000011101001111111000000000111110110100000001100000000000001010011011100100110000000101010111111111000011110010000111111000111111000100011011111000";
W(28)<="0000111110111001111010110001011001110101100000000011001010110111010100001011111010110100000000000000001011001011011010100010110010101110010010000011011000111110011000100010001110010111000000100001110001110100010000011110101011001110000010100101011111001111011001000100001001100001110000000000000000001111110100101111001000100001111010011001010001001000000100110100000100000000000000001001010110111110011001001101101110111011111001000001000000001010011101111110000010101110001110011000001001110100111100000111000110001000000000001100001101000101100010010000101100010000110000001011100001111000000000100000001100101110110001110000010000110100111010011100100000100101011001011111000001000110000100101010110110101111001001100000100000100000110101100111001001010110000000001111100000001011";
W(29)<="0010000000001100000001001001111011111111110000100001100010000001110001111111100001010000000000010001101111111111100000000110011101010111111000000001100001101110111111110000001100001101111111111101000011010110011001111111100000001110100100000001111110010000111101001000000001111110100011100011000000000001111010011000010101110000000011101000001000001111100000001110010000100011111111100000111111000001110111111111100000101110000111111111111110000011111100000011111010110000101011111000000011011110110010110111111100000000111101011111111111011101111010111111100101111001001111001101001010011111001110111101100000111100011100000011101111001110111011110110110111111011111111011101111000000000000111110110001110011000000000000001011101010001000100001000010110011001111000000100110010111011";
W(30)<="0111101001101010011001101010101110000000001001000100000110111001011000010110000000101001000010100000001010010001110010000000001010000000111011111101100000000000011011010001011111011100000011011111010000100001101100000000111101110000000000101011000000001011100000111000011001011000100111001000001100110000110000110100000001100001100001111111010000001100011011001101001110000010000000000110010101011111101110000010001111011101111010001000100001100011011001100000000100000100001110111000000000000000111010001000100100010000000001100001100001000000100000001100010110100000000000000010101001000100101000000100000001111010011000000000000101111110000110111100100001111111000100000010010111011011111101110000000100111001111111100110000011001111010001110110011000011110011100111110000011111011";
W(31)<="1011100100000000001001111110111100000000000000000000001101100000000000000000000010110100000000010110001000000001110000110000001000010000000000100111110110000000000010001010011000100000000000001001001100100111000000000001100000000000000000000000011110001100000000011110000111111010111010100111111100111011000111111111111111010011101000000110100110111101111111111101111100111111111111111111110111110111111111111111110000111110001000011001111101000001000001001011000011000000001010000111111100000000000000011000001011100000000000110101010011111100000001101000110001001110100000000001110010000011111111000000000111100000001111001111110001100100111101000111111101100010000001111000001010000000000000000111101000000001000000000001010100010000000110000000000111101000000010101100111001001000";
W(32)<="0101000101001100000000000111011000110110010101111100101101111111010101000000000001011011111111111001001100000100001111111111011110001000110100111010000000111101111011110011000011011111000010001110010000011010110100000110111111000011111111011110000010001000000001010011111100000101100001001111111111111010011010101000101111111111111101011011110000110111111111110110000111111011111110111111111000011111101111111111111000000001111111111011111001100000000111111111000111111110000100000111111000000000011000010000001111110000000000010001100000001011111000000011100110000000111111100011001111010000001010111111111111111010011000000010111111111111111001000011101111111111111111101010001111111101111111011111011011110110000001011100111101010011111000000000011011000001010110011000011000000111";
W(33)<="1101010100000100110110101010100110100000000000000010001000110110000000000000000011110110100111100000000011100100000000011111101101101110010010110000111101100011111111001011000011111100110111111000001100000101010110001001001110111000000000100000000000111011100000000111110000000010001100000000011111100000001010110000000011101011001001001100000000011110100110000000110000000001111100000001000101100000001111110000011100110110000000101111000000100100011111000001111000000010001101110000000111101000000001010110000101111110000000000001100000000000000000000000000100000001100000000000000000010001110100000000000000000001100111100100001010000000001110001100000000000110010000010110000000000000000011110000001000000000000000000111101100011101010101000011011110000000100101011110110001011001";
W(34)<="1101111111101111000010010100011011111111111111111110000000011111111101010111101110011001111111110100000011100111001111001011100111000000001110110001001111110111101000001010000000001111000000101000011000000001011000001100111111000000000000000000000011001100000000000011101110000111100000000000111110110000011000000000001111110100100101111000000011111111100000011010000000111111111100000101111000000111111111100000101111110000111111111100000011111011000001111111110111111111100010000111111110011111111010001000011111100111111111111100100001101100111000011111101001001100001110111111100110100010011011110111100000000010101110111010010110000000100011001111111000000000000000110010110000000000000000010111110100000000000000000000011100010000000000000000001111010010110010001000110011001011";
W(35)<="0010010101110000000001001100101000000000001111100001011011111110000001001000001111110111000010100000000000000011111000000111000001001110000111111000011100000001000000001011000000110100111100000000001100000101111111100000010100100000011101111111100000111010000001101111100001000011101000000011011001000010001100010000011001100110001000110000000000001111111101000001010000000001110101111110010100000000000001100011010000000100000000001111000000001000111111000000111100000000000011111111100111110000000100001111110111111111000000000000001101011111111000000000001000111111101101010000000000111011110000000000000000011100000111000000000000000010110110101010000000100000010100110100001110000000000000101001111011111100100000000110101000111111010011000010001001101011110101110100110011001010";
W(36)<="0110001000000100110110110001111000111110011111001001110101100111101111111111111111010110000000111111111111111000011000000000001101111111110011000000000011000110011111111000000011110111111111111011010110111101011111111111101111111011111111111111111111110011111111111000000010111111011111111111000000001111111001111111111001111110011111111111111101010011111110011111011110100100111111100000100100110000001101111000000010000000000000110110000000000111000000000000110000000000111011100000000010000000001011111110000000000000000011111110011000000000010101110111101011100000001010111011011110101110000101100110111111111110010100001001000011111101111100111110001111111111111111010111111111111111111111111110100111111111111111111000110000001111111111111111011101101110100011101111111111010101";
W(37)<="0100111000110100001000101101010000000000000000000001010101100000000000000000000001010111000000000000000100000010011111110000000110111111001101111111111110111111101111000111111111111101111010000101000111111111110111101110010011011111111111111110101100001011111111111111111110100000111111011111011111111110000111110111111101111111111000001111110010000001111111100001011110011001000011101110000000011010000000001010000001010001111001100000000100001000000011101000000000000000000000000101011000000000001001000000001100000000010010100101000001000000011011000010011100000010010000000000101001000000000000001001000010000011000110001000111100010001000010001101000000000000000000011111111110110110111000011011100001101011111111111110011001101011101100111111010001001000000101100111101111001001";
W(38)<="0010000000000000000000001101010010010110000110000000111011000001111010000100000000111100111111111111001000000001011111111111111111100000000001101111111111111111111000010100111111111111111111100011000011111110110000011110000000001101011000000010111000010001110100000000010000000100000100010000001111000001001110010000000001110000000000101000000000000110000000000011110000000000111001000000000111111101000010001011011000001111111010000101001011100101111111010000011101110010000001111111110001111101011001010111110000000010101011000001111110111101001011011100000010011110111111111101110000011011111111111011111000000000111001011111111111111000001101110100000011111111000011101100111000000000000000000011010001011000000000010000101110011000001110001001101010010010111000110110000110001101";
W(39)<="0101001001111111111111110110100000000000000000000010001101100000000000000000000011001110000000000011000000011001011000000001100000000001000010100000100100000000000000010110001000000000000000011101100000000001000000010001111101111000000001100000100101110111101111111110001011110010011111111111111001001101001101111111111111100101100110000111100001111110111111111110111110011111111111100011101111100011111010011101111001110110000000011011110100001100111000001011101111111101111111111111111111011111000111001011111111100000000010110110001111111000000001111110111011111100000000000010111111110111100000000000010111110000001111001111110111000010100111100000001000000000001000001000000000000000000000001000010000000001000000000001101001000000000010000000000001110100100111100000001001110110";
W(40)<="1001101100111110100100010001100110001111101100000011111101110001111101110111011101001001001011011110100001001101101100111010110101110001011000111100011010110010110101111011110100010101110001110000001010010000000000001011011110011000111100110000000101011110011000000100111001011111000011001101000001011001101111110000001000010000001110100010011001000011001111001110001000001100000011001010110111011110100010001010001000101110000000100010101010010000110011001010011001001001011101111111000000000000000001101110001011110000001011111101001111100000010000001101101110010011111010100001001010000010111100000101101110111011100000000001010111110100111110011010001000000001010011000011100001100111100110110111101100011001110010010100001100111101001001000101101010011010101101100100011010110011";
W(41)<="1010100000000111101111110100001011001000111111000001000010100100000000111111110100000111111100101111111001111000111111111111111011101111100101101111111111111011011111000110111111101111111111111100101001111101111111111111101111010110011111111011111110110100000111111001000011111111101000001100000000000111110100110110110000000111111110010111101100000000011111110000011011110100000001011010000000100010000000001100000001101000000100000000100000000010100000000000000000000000001010000001011000000000000001000010100111111000000000000100011011001011111100000001011111110111011111111100001111100111111111111111111110001110010110101101001111011011001000100011111100111111111110110011100111111111111111101100000111000111111111111110111011111111111100111011111000101000110000100011010111110010";
W(42)<="1010101110011000001111110010011110000000000000000000000011100000000000000000000000010111011111111101101000000010111110111111111101111100000001110011111011101111111111101111110111111111111111001110111111110111111111111111011011111111011111111111001100111011111001101111111110110011111111011000111111111011101111110010010111111110111110001110001000111111100000000000111001000011111110000000000011111101110111110010000000011111101101001100000000000010001111101000010001000011001000000000000000010110010100100000000000000100001010000010110000000000000000001001011110000010000000000001000000101000000000000010000000000000100111111111000000000001011000011111110001100001100001010011111111111111111111100111110111111111111111111111100011011111110111111111111011101111100100100000001100011111";
W(43)<="1110100000000000000000101100000000000000000000000000001010101100000000000000000011101000000011010001111000000010100000011111111101110111001110001100111111101100101100010000011001101111101100000011000000000111110101111000001010000010000010111100000000111000000011011111101000000011000010010100011111110000001100001010100111111011100000100001110110001111101111001110000111100010111011001110111100011110100011111111110000010001100001111111111111000001111110000000011111111000001101110000000000111111100000010111101000000000111110000000111111100000000011111000000100111000000000001101100001010011100000000000010010000110101111111111010100100000011001111111100000000001010010001011111111110010011111101001110111111111111111111111101111100111110000111011111101001100010110000010010101101010";
W(44)<="0111111111111111101001010110001001111111111111111111111000010011111111111111111100011100000000101100110000100011100000001010001110000000001110110000011010011000000000000010000000111011100000000000100000000100111110000000010010000000000001110000000011011000000001011111110000000111000000111001110011100000110100000111110111000111100001011000011111111100110011000001000011100100110001000100000000000011111101000110001111110000000101100111101111111111000001100100011101011011111010000100000011111001111111101100000000011111111111111110000000000001111111011011111000000000000111110000001111100000000000010000001111011101110000000000000010100111111000000001111000111101111111000010111111111111111111111110111111111111111111111110011011111111110111111111111111101010110010100011011010100111";
W(45)<="1101000001111100000000011011111000010100000100011101110101011111010101111111100001101011111101101000010111000000110111111100000000000000000110111001100100000000000000100010000111111111000000000111101000000111111110000000001100000000000101100000000000001000000110111111110000000001000000011101111111110000000100000001101111011111100000100000010111111111111110001110000000111111111111111111111000000010111111111111111110010000000111111111111111110000000000001100000111111010000000000000000000000011000000010000000000000000001010000001000000000000101000000011000001000000010000000000000000010100110000000000000001110111000111110100000000010101001011011111101000000000111100101111111111101100111111010010001001100001000001110011110000010100001110000001101110100001110001110000110011101111";
W(46)<="1011111111111111111111110000011111111111111011111110101101110111111111111111111111001000000000110111110011111000110000000111011010111111100101000000101110111011111011010100000000000001101101111101100000000000001110010111101101000010000000010101111111100110011011100000010000010110111111101111000000100111011011001111110100000111101101011101111111000000010010100111011110111100000000000000011010111100000000000000000001101001110010110000000000001110000011111111100000000001111000001111111111111100001111110000011111111111010110111100000001011111111111111111101100000011011101111111111111110000001010010111111111111101000000001001111111111111111110000000111010111111101111001100000000001001100000110010111101100000000000001011000011010100001100011100011011110000000000110100110010110110";
W(47)<="0001000000001000000000010111111011111100000000000001001000000000100000001110111111101000000000111111111110011011110100000001111111110011111111000000001111111110010011011100000001000010111011111011100000000010101011111111101100000001011100000011111011110000010011111000000111111110000001101111000000011111101010011100011000000000011111100001111000000001110000110110000111000000001110000000111100001000000101111000000010000111000000101111110000000001111110000111011111010000000011111111110101111111000011111111111110100100111100000000011111111101000110101100000111111100011011010000000000101111110100101111000111110011011110110111011011011110100111111100000010111101111111111101100000100001000001101111101000011110000000000110011010000110000000110101001010011001101110000100111100110100";
W(48)<="1000100100111110011110011100011001111000011101000010011110001101101110111111111101100110011101100111111111111000011100000110101111111111110001001111101101010010001110111000001101101111000110011111000000110111010000011111101110000111111000000000011111101000011111110000000000011110000001111000000000000001111000000111100000010000000011110000001110010011100000001101010000011000110100100001100111000000010101111000000110000110000000010111000000011101010000000000000000000000110011100000000000000000111111001110000000000010000000011101111100001111110010100011101111111111111111000000000110101111111110101111110000011100011111001110000101000010100011111111111111001001111111011101111111111000000001010110111011111111111100011100010000001111111001111011111010000000101010110111111001001110";
W(49)<="0010000000001000000000001011000110011111111110001001110100000001111101001000000001111000010111111000011100000001100011111111111110100000001101001111011111111000001000101100111101101111110111100001110000011010111111110010011000000100011010111111100001010000000000000011111111100001000111010000000111110110000000011000000000011111010110000000100000000001011100100011000111100000001111000000000100001110000110111111110000100001111000100111111111000011111111100000001111111100010011111100000000111111110011000111101010000111111110000100111111100101111010110000000010111000011111100101000000001011100110111101101000000010011011111111110010000000001010111111010111100000000000101111111010001110000000000100101101111111111111101110100111011111111110111111110011010101111110011111110010101110";

	TO_INTEGER_i:
	for i in 0 to N_INPUTS generate  
	begin
		INTEGER_INPUT(i) <= (to_integer(unsigned(INPUT(i)))); 
	end generate;
	
	W_DOT_INPUT_i:
	for i in 0 to N_OUTPUTS generate  
	begin
		INTEGER_W_DOT_INPUT_j:
		for j in 0 to N_INPUTS generate  
		begin
			INTEGER_W_DOT_INPUT(i)(j) <= -INTEGER_INPUT(j) when W(i)(j) = '0' else INTEGER_INPUT(j);  
		end generate;
		
		W_DOT_INPUT(i) <= f_sum(INTEGER_W_DOT_INPUT(i));
	end generate;
	
	RELU_i:
	for i in 0 to N_OUTPUTS generate  
	begin
		RELU(i) <= W_DOT_INPUT(i) when W_DOT_INPUT(i) > 0 else 0;
	end generate;

	NORMALIZED_BATCH_i:
	for i in 0 to N_OUTPUTS generate
	begin
		NORMALIZED_BATCH(i) <= GAMMA(i) * (RELU(i) - MEAN(i)) / STD_DEV(i) + BETA(i);
	end generate;
	
	
	OUTPUT_i:
	for i in 0 to N_OUTPUTS generate  
	begin
		OUTPUT(i) <= '1' when (NORMALIZED_BATCH(i) > 0) else '0';
	end generate;
	
end layer;
